// Universidad del Valle de Guatemala
// Valerie Valdez

//                    Electrónica digital
//                     Laboratorio No. 10
//                       Ejercicio No. 2


// Testbench
module testbench();
  input wire;
